library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
    port(
        clk: in std_logic;
        address: in unsigned(6 downto 0);
        data : out unsigned(14 downto 0)
    );
end entity;

architecture a_rom of rom is
    type rom_array_type is array (0 to 127) of unsigned(14 downto 0);

    signal rom_memory : rom_array_type := (
       -- ============================================================
        -- FASE 1: INICIALIZAÇÃO
        -- ============================================================
        0  => "0001" & "1000" & "0000000", -- 0: CLR R8
        1  => "0101" & "1000" & "0100000", -- 1: ADDI R8, 32
        
        2  => "0001" & "0001" & "0000000", -- 2: CLR R1
        3  => "0101" & "0001" & "0000001", -- 3: ADDI R1, 1

        -- LOOP INIT (Addr 4)
        -- SW R1, R1 -> Endereço R1 (Rx), Dado R1 (Ry). OK!
        4  => "1010" & "0001" & "0001" & "000", 
        5  => "0101" & "0001" & "0000001", 
        6  => "0010" & "0111" & "0001" & "000", 
        7  => "0100" & "0111" & "1000" & "000", 
        
        8  => "0111" & "0000" & "1111100", 
        9  => "0000" & "0000" & "0000000", 

        -- ============================================================
        -- FASE 2: FILTROS
        -- ============================================================
        10 => "0001" & "0000" & "0000000", -- 10: CLR R0

        -- --- FILTRO DO 2 ---
        11 => "0001" & "0010" & "0000000", -- 11: CLR R2
        12 => "0101" & "0010" & "0000100", -- 12: ADDI R2, 4

        -- LOOP CHECK 2 (Addr 13)
        13 => "0010" & "0111" & "0010" & "000", 
        14 => "0100" & "0111" & "1000" & "000", 
        
        15 => "0111" & "0000" & "0000100", 
        16 => "0000" & "0000" & "0000000", 
        
        17 => "0110" & "0000" & "0010111", 
        18 => "0000" & "0000" & "0000000", 

        -- APAGAR 2 (Addr 19)
        -- CORRIGIDO: SW R2(Addr), R0(Data)
        -- Antes: "1010" & "0000" & "0010" -> Agora: "1010" & "0010" & "0000"
        19 => "1010" & "0010" & "0000" & "000", 
        
        20 => "0101" & "0010" & "0000010", 
        
        21 => "0110" & "0000" & "0001101", 
        22 => "0000" & "0000" & "0000000", 

        -- --- FILTRO DO 3 --- (Addr 23)
        23 => "0001" & "0010" & "0000000", 
        24 => "0101" & "0010" & "0000110", 

        -- LOOP CHECK 3 (Addr 25)
        25 => "0010" & "0111" & "0010" & "000", 
        26 => "0100" & "0111" & "1000" & "000", 
        
        27 => "0111" & "0000" & "0000100", 
        28 => "0000" & "0000" & "0000000", 
        
        29 => "0110" & "0000" & "0100011", 
        30 => "0000" & "0000" & "0000000", 

        -- APAGAR 3 (Addr 31)
        -- CORRIGIDO: SW R2(Addr), R0(Data)
        31 => "1010" & "0010" & "0000" & "000", 
        
        32 => "0101" & "0010" & "0000011", 
        
        33 => "0110" & "0000" & "0011001", 
        34 => "0000" & "0000" & "0000000", 

        -- --- FILTRO DO 5 --- (Addr 35)
        35 => "0001" & "0010" & "0000000", 
        36 => "0101" & "0010" & "0001010", 

        -- LOOP CHECK 5 (Addr 37)
        37 => "0010" & "0111" & "0010" & "000", 
        38 => "0100" & "0111" & "1000" & "000", 
        
        39 => "0111" & "0000" & "0000100", 
        40 => "0000" & "0000" & "0000000", 
        
        41 => "0110" & "0000" & "0101111", 
        42 => "0000" & "0000" & "0000000", 

        -- APAGAR 5 (Addr 43)
        -- CORRIGIDO: SW R2(Addr), R0(Data)
        43 => "1010" & "0010" & "0000" & "000", 
        
        44 => "0101" & "0010" & "0000101", 
        
        45 => "0110" & "0000" & "0100101", 
        46 => "0000" & "0000" & "0000000", 

        -- ============================================================
        -- FASE 3: LEITURA E DISPLAY
        -- ============================================================
        47 => "0001" & "0001" & "0000000", 
        48 => "0101" & "0001" & "0000010", 

        -- LOOP LEITURA (Addr 49)
        -- LW R4, (R1) -> Op(1001) | Dest R4(Rx) | Addr R1(Ry).
        -- Rx=0100, Ry=0001. ESTA CORRETO COM A NOVA ARQUITETURA!
        49 => "1001" & "0100" & "0001" & "000", 
        
        50 => "0000" & "0000" & "0000000", 
        
        51 => "0010" & "0110" & "0100" & "000", 
        
        52 => "0101" & "0001" & "0000001", 
        53 => "0010" & "0111" & "0001" & "000", 
        54 => "0100" & "0111" & "1000" & "000", 

        55 => "0111" & "0000" & "1111010", 
        56 => "0000" & "0000" & "0000000", 

        57 => "0110" & "0000" & "0111001", 
        58 => "0000" & "0000" & "0000000", 
        
        others => (others => '0')
    );
begin
    process(clk)
    begin
        if rising_edge(clk) then
            data <= rom_memory(to_integer(address));
        end if;
    end process;
end architecture a_rom;